----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:33:48 04/23/2014 
-- Design Name: 
-- Module Name:    Four_min_struct - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
LIBRARY ieee ;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
 
ENTITY four_min IS
   PORT(
      clk         : IN     std_logic  ;
      dat_in0     : IN     std_logic_vector (7 DOWNTO 0) ;
      dat_in1     : IN     std_logic_vector (7 DOWNTO 0) ;
      dat_in2     : IN     std_logic_vector (7 DOWNTO 0) ;
      dat_in3     : IN     std_logic_vector (7 DOWNTO 0) ;
      en          : IN     std_logic  ;
      dat_out     : OUT    std_logic_vector (7 DOWNTO 0) ;
      dat_out_pos : OUT    std_logic_vector (1 DOWNTO 0)
   );
 
-- Declarations
 
END four_min ;
 
-- renoir interface_end
--
-- VHDL Architecture Comparer.four_min.struct
--
-- Created:
--          by - sweather.UNKNOWN (SWMOBL)
--          at - 15:16:33 05/09/2001
--
-- Generated by Mentor Graphics' Renoir(TM) 2000.3 (Build 2)
--
LIBRARY ieee ;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
 
LIBRARY Comparer;
 
ARCHITECTURE struct OF four_min IS
 
   -- Architecture declarations
 
   -- Internal signal declarations
   SIGNAL dbus10 : std_logic_vector(7 DOWNTO 0);
   SIGNAL dbus12 : std_logic_vector(7 DOWNTO 0);
   SIGNAL dbus13 : std_logic_vector(1 DOWNTO 0);
   SIGNAL dbus14 : std_logic_vector(7 DOWNTO 0);
   SIGNAL dbus15 : std_logic_vector(1 DOWNTO 0);
   SIGNAL dbus4  : std_logic_vector(7 DOWNTO 0);
   SIGNAL dbus6  : std_logic_vector(7 DOWNTO 0);
   SIGNAL dbus8  : std_logic_vector(7 DOWNTO 0);
 
   -- Component Declarations
   COMPONENT Compare0
   PORT (
      dbus4  : IN     std_logic_vector (7 DOWNTO 0);
      dbus6  : IN     std_logic_vector (7 DOWNTO 0);
      dbus12 : OUT    std_logic_vector (7 DOWNTO 0);
      dbus13 : OUT    std_logic_vector (1 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT Compare1
   PORT (
      dbus10 : IN     std_logic_vector (7 DOWNTO 0);
      dbus8  : IN     std_logic_vector (7 DOWNTO 0);
      dbus14 : OUT    std_logic_vector (7 DOWNTO 0);
      dbus15 : OUT    std_logic_vector (1 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT Compare3
   PORT (
      dbus12      : IN     std_logic_vector (7 DOWNTO 0);
      dbus13      : IN     std_logic_vector (1 DOWNTO 0);
      dbus14      : IN     std_logic_vector (7 DOWNTO 0);
      dbus15      : IN     std_logic_vector (1 DOWNTO 0);
      dat_out     : OUT    std_logic_vector (7 DOWNTO 0);
      dat_out_pos : OUT    std_logic_vector (1 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT latch0
   PORT (
      clk     : IN     std_logic ;
      dat_in0 : IN     std_logic_vector (7 DOWNTO 0);
      en      : IN     std_logic ;
      dbus4   : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT latch1
   PORT (
      clk     : IN     std_logic ;
      dat_in1 : IN     std_logic_vector (7 DOWNTO 0);
      en      : IN     std_logic ;
      dbus6   : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT latch2
   PORT (
      clk     : IN     std_logic ;
      dat_in2 : IN     std_logic_vector (7 DOWNTO 0);
      en      : IN     std_logic ;
      dbus8   : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT latch3
   PORT (
      clk     : IN     std_logic ;
      dat_in3 : IN     std_logic_vector (7 DOWNTO 0);
      en      : IN     std_logic ;
      dbus10  : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;
 
   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Compare0 USE ENTITY Comparer.Compare0;
   FOR ALL : Compare1 USE ENTITY Comparer.Compare1;
   FOR ALL : Compare3 USE ENTITY Comparer.Compare3;
   FOR ALL : latch0 USE ENTITY Comparer.latch0;
   FOR ALL : latch1 USE ENTITY Comparer.latch1;
   FOR ALL : latch2 USE ENTITY Comparer.latch2;
   FOR ALL : latch3 USE ENTITY Comparer.latch3;
   -- pragma synthesis_on
 
BEGIN
   -- Instance port mappings.
   I4 : Compare0
      PORT MAP (
         dbus4  => dbus4,
         dbus6  => dbus6,
         dbus12 => dbus12,
         dbus13 => dbus13
      );
   I5 : Compare1
      PORT MAP (
         dbus10 => dbus10,
         dbus8  => dbus8,
         dbus14 => dbus14,
         dbus15 => dbus15
      );
   I6 : Compare3
      PORT MAP (
         dbus12      => dbus12,
         dbus13      => dbus13,
         dbus14      => dbus14,
         dbus15      => dbus15,
         dat_out     => dat_out,
         dat_out_pos => dat_out_pos
      );
   I0 : latch0
      PORT MAP (
         clk     => clk,
         dat_in0 => dat_in0,
         en      => en,
         dbus4   => dbus4
      );
   I1 : latch1
      PORT MAP (
         clk     => clk,
         dat_in1 => dat_in1,
         en      => en,
         dbus6   => dbus6
      );
   I2 : latch2
      PORT MAP (
         clk     => clk,
         dat_in2 => dat_in2,
         en      => en,
         dbus8   => dbus8
      );
   I3 : latch3
      PORT MAP (
         clk     => clk,
         dat_in3 => dat_in3,
         en      => en,
         dbus10  => dbus10
      );
 
END struct;

