INFO:HDLCompiler:1061 - Parsing VHDL file "/home/cccitron/mastersThesis/makestuff/libs/libfpgalink-20120621/hdl/fx2/vhdl/sad_simple_reg_3x3/top_level/sad_wrapper.vhd" into library work
INFO:ProjectMgmt - Parsing design hierarchy completed successfully.
INFO:HDLCompiler:1061 - Parsing VHDL file "/home/cccitron/mastersThesis/makestuff/libs/libfpgalink-20120621/hdl/fx2/vhdl/sad_simple_reg_3x3/top_level/sad_wrapper.vhd" into library work
INFO:ProjectMgmt - Parsing design hierarchy completed successfully.
